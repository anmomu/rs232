module top ();


endmodule
